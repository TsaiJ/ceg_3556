ROM_1_port_lab2_inst : ROM_1_port_lab2 PORT MAP (
		address	 => address_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
